`timescale 1ns / 1ps

module alu_control(
  input [3:0] funct3,
  input [6:0] funct7,
  input [6:0] opcode,
  output [3:0] alu_op
);


endmodule