`define ADD 4'h0
`define SLL 4'h1
`define SLT 4'h2
`define SLTU 4'h3
`define XOR 4'h4
`define SRL 4'h5
`define OR  4'h6
`define AND 4'h7

`define SUB 4'hA
`define SRA 4'hD

`define ALU_OP_MEM  2'b00
`define ALU_OP_BEQ  2'b01
`define ALU_OP_MATH 2'b10


