`timescale 1ns / 1ps

module cpu_tb();



endmodule