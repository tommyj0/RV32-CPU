`define ADD 4'h0
`define SUB 4'h1
`define AND 4'h2
`define OR  4'h3
`define XOR 4'h4
`define SLL 4'h5
`define SRL 4'h6
`define SRA 4'h7


`define MUL 4'hD
`define DIV 4'hE
`define REM 4'hF
