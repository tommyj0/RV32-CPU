`define	QUAD_MASK		32'hc0000000
`define	ROM_BASE_ADDR		32'h0
`define	RAM_BASE_ADDR		32'h40000000
`define	EXT_BASE_ADDR		32'h80000000
`define	IO_BASE_ADDR		32'hc0000000
`define	VGA_ADDR		32'hc0000000
