`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
//
// MODULE: CPU
//
////////////////////////////////////////////////////////////////////////////////



module cpu(

    );
endmodule